digraph finite_state_machine {
	rankdir=LR;
	size="8,5"
	node [shape = circle];
	start -> price-pos [ label = "0.1983050847" ];
	start -> servic-pos [ label = "0.0618644068" ];
	start -> picture-pos [ label = "0.0779661017" ];
	start -> quality-pos [ label = "0.0983050847" ];
	start -> price-neg [ label = "0.1271186441" ];
	start -> quality-neg [ label = "0.0584745763" ];
	screen-pos -> price-pos [ label = "0.5033557047" ];
	screen-pos -> sound-pos [ label = "0.1006711409" ];
	screen-pos -> quality-pos [ label = "0.0648769575" ];
	screen-pos -> app-pos [ label = "0.0648769575" ];
	screen-pos -> screen-neg [ label = "0.0760626398" ];
	price-pos -> price-pos [ label = "0.0541436464" ];
	price-pos -> sound-pos [ label = "0.5546961326" ];
	price-pos -> picture-pos [ label = "0.0740331492" ];
	price-pos -> quality-pos [ label = "0.070718232" ];
	price-pos -> screen-neg [ label = "0.0651933702" ];
	sound-pos -> sound-pos [ label = "0.0523690773" ];
	sound-pos -> servic-pos [ label = "0.5436408978" ];
	sound-pos -> quality-pos [ label = "0.0673316708" ];
	sound-pos -> screen-neg [ label = "0.0972568579" ];
	servic-pos -> sound-pos [ label = "0.0833333333" ];
	servic-pos -> picture-pos [ label = "0.6914893617" ];
	picture-pos -> price-pos [ label = "0.0775444265" ];
	picture-pos -> sound-pos [ label = "0.0694668821" ];
	picture-pos -> servic-pos [ label = "0.0533117932" ];
	picture-pos -> quality-pos [ label = "0.5201938611" ];
	picture-pos -> screen-neg [ label = "0.0743134087" ];
	quality-pos -> sound-pos [ label = "0.0727272727" ];
	quality-pos -> picture-pos [ label = "0.0613636364" ];
	quality-pos -> quality-pos [ label = "0.0704545455" ];
	quality-pos -> app-pos [ label = "0.5136363636" ];
	app-pos -> servic-pos [ label = "0.0555555556" ];
	app-pos -> picture-pos [ label = "0.0555555556" ];
	app-pos -> quality-pos [ label = "0.0740740741" ];
	app-pos -> app-pos [ label = "0.0740740741" ];
	app-pos -> connection-pos [ label = "0.462962963" ];
	app-pos -> screen-neg [ label = "0.0648148148" ];
	connection-pos -> price-pos [ label = "0.0540935673" ];
	connection-pos -> screen-neg [ label = "0.6286549708" ];
	screen-neg -> price-neg [ label = "0.5426829268" ];
	screen-neg -> sound-neg [ label = "0.0884146341" ];
	screen-neg -> picture-neg [ label = "0.1082317073" ];
	screen-neg -> quality-neg [ label = "0.0579268293" ];
	price-neg -> price-neg [ label = "0.0602678571" ];
	price-neg -> sound-neg [ label = "0.6104910714" ];
	price-neg -> picture-neg [ label = "0.0993303571" ];
	price-neg -> quality-neg [ label = "0.0502232143" ];
	sound-neg -> price-neg [ label = "0.0619047619" ];
	sound-neg -> sound-neg [ label = "0.0619047619" ];
	sound-neg -> servic-neg [ label = "0.5666666667" ];
	sound-neg -> picture-neg [ label = "0.0619047619" ];
	sound-neg -> quality-neg [ label = "0.0547619048" ];
	servic-neg -> sound-neg [ label = "0.0898989899" ];
	servic-neg -> picture-neg [ label = "0.7101010101" ];
	picture-neg -> price-neg [ label = "0.0603085554" ];
	picture-neg -> sound-neg [ label = "0.0532959327" ];
	picture-neg -> servic-neg [ label = "0.0532959327" ];
	picture-neg -> quality-neg [ label = "0.6100981767" ];
	quality-neg -> price-neg [ label = "0.0780141844" ];
	quality-neg -> sound-neg [ label = "0.0945626478" ];
	quality-neg -> picture-neg [ label = "0.0969267139" ];
	quality-neg -> quality-neg [ label = "0.0638297872" ];
	quality-neg -> app-neg [ label = "0.4846335697" ];
	app-neg -> connection-neg [ label = "0.685560054" ];
	connection-neg -> picture-neg [ label = "0.0524553571" ];
	connection-neg -> connection-neg [ label = "0.0636160714" ];
}
