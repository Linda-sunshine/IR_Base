digraph finite_state_machine {
	rankdir=LR;
	size="8,5"
	node [shape = circle];
	start -> zoom-pos [ label = "0.0917797287" ];
	start -> picture-pos [ label = "0.0662410215" ];
	start -> price-pos [ label = "0.1476456504" ];
	start -> Instruction-pos [ label = "0.0582601756" ];
	start -> zoom-neg [ label = "0.0526735834" ];
	start -> picture-neg [ label = "0.0734237829" ];
	start -> price-neg [ label = "0.0845969673" ];
	battery-pos -> screen-pos [ label = "0.4599406528" ];
	battery-pos -> zoom-pos [ label = "0.056379822" ];
	battery-pos -> price-pos [ label = "0.0534124629" ];
	battery-pos -> Instruction-pos [ label = "0.059347181" ];
	screen-pos -> screen-pos [ label = "0.0555555556" ];
	screen-pos -> viewfinder-pos [ label = "0.2777777778" ];
	screen-pos -> len-pos [ label = "0.0714285714" ];
	screen-pos -> picture-pos [ label = "0.0634920635" ];
	screen-pos -> price-pos [ label = "0.0873015873" ];
	screen-pos -> Instruction-pos [ label = "0.0714285714" ];
	screen-pos -> video-pos [ label = "0.0555555556" ];
	viewfinder-pos -> record-pos [ label = "0.3376623377" ];
	viewfinder-pos -> len-pos [ label = "0.0584415584" ];
	viewfinder-pos -> picture-pos [ label = "0.0649350649" ];
	viewfinder-pos -> price-pos [ label = "0.0909090909" ];
	viewfinder-pos -> Instruction-pos [ label = "0.0714285714" ];
	viewfinder-pos -> video-pos [ label = "0.0584415584" ];
	record-pos -> screen-pos [ label = "0.0714285714" ];
	record-pos -> mode-pos [ label = "0.3979591837" ];
	record-pos -> shutter-pos [ label = "0.0714285714" ];
	record-pos -> price-pos [ label = "0.0816326531" ];
	record-pos -> Instruction-pos [ label = "0.0714285714" ];
	record-pos -> video-pos [ label = "0.0612244898" ];
	mode-pos -> shutter-pos [ label = "0.4393638171" ];
	mode-pos -> len-pos [ label = "0.0536779324" ];
	mode-pos -> picture-pos [ label = "0.0675944334" ];
	mode-pos -> price-pos [ label = "0.0715705765" ];
	shutter-pos -> shutter-pos [ label = "0.0762711864" ];
	shutter-pos -> memori-pos [ label = "0.3728813559" ];
	shutter-pos -> picture-pos [ label = "0.0847457627" ];
	shutter-pos -> price-pos [ label = "0.1228813559" ];
	memori-pos -> screen-pos [ label = "0.0765957447" ];
	memori-pos -> shutter-pos [ label = "0.0723404255" ];
	memori-pos -> zoom-pos [ label = "0.3829787234" ];
	memori-pos -> Instruction-pos [ label = "0.0638297872" ];
	memori-pos -> video-pos [ label = "0.0510638298" ];
	memori-pos -> battery-neg [ label = "0.0553191489" ];
	zoom-pos -> len-pos [ label = "0.403887689" ];
	zoom-pos -> picture-pos [ label = "0.0583153348" ];
	zoom-pos -> price-pos [ label = "0.090712743" ];
	zoom-pos -> Instruction-pos [ label = "0.0691144708" ];
	len-pos -> shutter-pos [ label = "0.0684210526" ];
	len-pos -> picture-pos [ label = "0.5333333333" ];
	len-pos -> price-pos [ label = "0.0666666667" ];
	len-pos -> video-pos [ label = "0.050877193" ];
	picture-pos -> shutter-pos [ label = "0.0653594771" ];
	picture-pos -> picture-pos [ label = "0.0640522876" ];
	picture-pos -> price-pos [ label = "0.4836601307" ];
	price-pos -> len-pos [ label = "0.0751879699" ];
	price-pos -> price-pos [ label = "0.0721804511" ];
	price-pos -> Instruction-pos [ label = "0.4766917293" ];
	price-pos -> video-pos [ label = "0.0601503759" ];
	Instruction-pos -> shutter-pos [ label = "0.0742574257" ];
	Instruction-pos -> picture-pos [ label = "0.0544554455" ];
	Instruction-pos -> price-pos [ label = "0.0668316832" ];
	Instruction-pos -> Instruction-pos [ label = "0.0792079208" ];
	Instruction-pos -> video-pos [ label = "0.3787128713" ];
	video-pos -> price-pos [ label = "0.0744680851" ];
	video-pos -> Instruction-pos [ label = "0.0567375887" ];
	video-pos -> battery-neg [ label = "0.4574468085" ];
	battery-neg -> screen-neg [ label = "0.4978991597" ];
	battery-neg -> mode-neg [ label = "0.0567226891" ];
	battery-neg -> Instruction-neg [ label = "0.1323529412" ];
	screen-neg -> viewfinder-neg [ label = "0.3045977011" ];
	screen-neg -> record-neg [ label = "0.0574712644" ];
	screen-neg -> shutter-neg [ label = "0.1091954023" ];
	screen-neg -> zoom-neg [ label = "0.0517241379" ];
	screen-neg -> price-neg [ label = "0.091954023" ];
	screen-neg -> Instruction-neg [ label = "0.0747126437" ];
	viewfinder-neg -> record-neg [ label = "0.3575418994" ];
	viewfinder-neg -> shutter-neg [ label = "0.094972067" ];
	viewfinder-neg -> len-neg [ label = "0.0726256983" ];
	viewfinder-neg -> price-neg [ label = "0.061452514" ];
	viewfinder-neg -> Instruction-neg [ label = "0.0502793296" ];
	record-neg -> mode-neg [ label = "0.4720496894" ];
	record-neg -> Instruction-neg [ label = "0.1583850932" ];
	mode-neg -> shutter-neg [ label = "0.5238095238" ];
	mode-neg -> price-neg [ label = "0.0952380952" ];
	shutter-neg -> shutter-neg [ label = "0.0825688073" ];
	shutter-neg -> memori-neg [ label = "0.4403669725" ];
	shutter-neg -> price-neg [ label = "0.0733944954" ];
	shutter-neg -> Instruction-neg [ label = "0.0642201835" ];
	memori-neg -> mode-neg [ label = "0.0502645503" ];
	memori-neg -> zoom-neg [ label = "0.5608465608" ];
	memori-neg -> price-neg [ label = "0.0555555556" ];
	memori-neg -> Instruction-neg [ label = "0.0925925926" ];
	zoom-neg -> shutter-neg [ label = "0.0939086294" ];
	zoom-neg -> len-neg [ label = "0.4111675127" ];
	zoom-neg -> price-neg [ label = "0.1116751269" ];
	zoom-neg -> Instruction-neg [ label = "0.0659898477" ];
	len-neg -> screen-neg [ label = "0.0597484277" ];
	len-neg -> shutter-neg [ label = "0.0628930818" ];
	len-neg -> picture-neg [ label = "0.3962264151" ];
	len-neg -> price-neg [ label = "0.0534591195" ];
	len-neg -> Instruction-neg [ label = "0.072327044" ];
	picture-neg -> shutter-neg [ label = "0.0769230769" ];
	picture-neg -> price-neg [ label = "0.552238806" ];
	picture-neg -> Instruction-neg [ label = "0.05510907" ];
	price-neg -> screen-neg [ label = "0.0857946554" ];
	price-neg -> price-neg [ label = "0.0604781997" ];
	price-neg -> Instruction-neg [ label = "0.5203938115" ];
	Instruction-neg -> shutter-neg [ label = "0.0633484163" ];
	Instruction-neg -> zoom-neg [ label = "0.0542986425" ];
	Instruction-neg -> price-neg [ label = "0.0678733032" ];
	Instruction-neg -> Instruction-neg [ label = "0.0633484163" ];
	Instruction-neg -> video-neg [ label = "0.3981900452" ];
	video-neg -> price-neg [ label = "0.071197411" ];
	video-neg -> Instruction-neg [ label = "0.1067961165" ];
}
